typedef enum logic[3:0] { //alu_ops
  ADD = 4'b1000;
  SUB = 4'b1001;
  INC = 4'b0110;
} alu_op;