module Controls(
    input carry,
    input [3:0] instruct_in,
    
)
endmodule: Controls